/*
* Top level design of the FPGC4
*/
module FPGC4(
    input clk, nreset,

    //VGA for GM7123 module
    output vga_hs,
    output vga_vs,
    output wire [7:0] vga_r,
    output wire [7:0] vga_g,
    output wire [7:0] vga_b,
    output wire VGAclk,
    output blk
);


endmodule